

module and_gate( a, b, y);
  input a, b; // input ports
  output y;  // output ports
  
  assign y = a & b ; // (a and b )
  
endmodule // no semicolon